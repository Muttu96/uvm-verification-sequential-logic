package counter_pkg;

        import uvm_pkg::*;
        `include "uvm_macros.svh"

        `include "agent_config.sv"

        `include "counter_xtn.sv"

        `include "sequence.sv"
        `include "sequencer.sv"
        `include "monitor.sv"
        `include "driver.sv"
        `include "agent.sv"

        `include "scoreboard.sv"

        `include "env.sv"
        `include "test.sv"

endpackage
