package dff_pkg;

        import uvm_pkg::*;
        `include "uvm_macros.svh"

        `include "agent_config.sv"

        `include "dff_transaction.sv"

        `include "dff_sequence.sv"
        `include "dff_sequencer.sv"
        `include "dff_monitor.sv"
        `include "dff_driver.sv"
        `include "dff_agent.sv"

        `include "dff_scoreboard.sv"

        `include "dff_env.sv"
        `include "dff_test.sv"

endpackage
